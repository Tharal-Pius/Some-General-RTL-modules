`include "transmitter.svh"
`include "double_flop_synch.svh"
`include "bin_to_gray.svh"
`include "gray_to_bin.svh"