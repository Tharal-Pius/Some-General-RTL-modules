`include "transmitter.sv"
`include "double_flop_synch.sv"
`include "bin_to_gray.sv"
`include "gray_to_bin.sv"